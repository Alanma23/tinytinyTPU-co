`timescale 1ns / 1ps

module pe (
    input  logic        clk,
    input  logic        reset,
    input  logic        en_weight_pass,    // Pass in_psum through out_psum (always during load phase)
    input  logic        en_weight_capture, // Capture weight from in_psum (per-PE timing for diagonal)
    input  logic signed [7:0]  in_act,
    input  logic signed [15:0] in_psum,
    output logic signed [7:0]  out_act,
    output logic signed [15:0] out_psum
);

    logic signed [7:0] weight;

    always_ff @(posedge clk) begin
        if (reset) begin
            out_act <= 8'sd0;
            out_psum <= 16'sd0;
            weight <= 8'sd0;
        end
        else begin
            if (en_weight_pass) begin
                // Weight loading mode: pass psum through, reset activation
                out_psum <= in_psum;
                out_act <= 8'sd0;
                // Capture weight only when this PE's capture signal is active
                if (en_weight_capture) begin
                    weight <= $signed(in_psum[7:0]);
                end
            end
            else begin
                // Compute mode: MAC operation (signed multiplication)
                out_act <= in_act;
                out_psum <= ($signed(in_act) * $signed(weight)) + in_psum;
            end
        end
    end

endmodule

